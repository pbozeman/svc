`ifndef SVC_RV_SOC_SRAM_SV
`define SVC_RV_SOC_SRAM_SV

`include "svc.sv"

`include "svc_mem_sram.sv"
`include "svc_rv.sv"

//
// RISC-V SoC with SRAM memories
//
// Single-cycle RISC-V core with separate instruction and data SRAMs.
// Both memories have 0-cycle read latency (combinational reads).
//
module svc_rv_soc_sram #(
    parameter int XLEN        = 32,
    parameter int IMEM_AW     = 10,
    parameter int DMEM_AW     = 10,
    parameter int IF_ID_REG   = 0,
    parameter int ID_EX_REG   = 0,
    parameter int EX_MEM_REG  = 0,
    parameter int MEM_WB_REG  = 0,
    parameter int REGFILE_FWD = 1,

    // verilog_lint: waive explicit-parameter-storage-type
    parameter IMEM_INIT = ""
) (
    input logic clk,
    input logic rst_n,

    output logic ebreak
);
  //
  // Memory interface signals
  //
  logic [31:0] imem_addr;
  logic [31:0] imem_data;

  logic [31:0] dmem_addr;
  logic [31:0] dmem_rdata;
  logic [31:0] dmem_waddr;
  logic [31:0] dmem_wdata;
  logic [ 3:0] dmem_wstrb;
  logic        dmem_we;

  //
  // RISC-V core
  //
  svc_rv #(
      .XLEN       (XLEN),
      .IMEM_AW    (IMEM_AW),
      .DMEM_AW    (DMEM_AW),
      .IF_ID_REG  (IF_ID_REG),
      .ID_EX_REG  (ID_EX_REG),
      .EX_MEM_REG (EX_MEM_REG),
      .MEM_WB_REG (MEM_WB_REG),
      .REGFILE_FWD(REGFILE_FWD)
  ) cpu (
      .clk       (clk),
      .rst_n     (rst_n),
      .imem_addr (imem_addr),
      .imem_data (imem_data),
      .dmem_addr (dmem_addr),
      .dmem_rdata(dmem_rdata),
      .dmem_waddr(dmem_waddr),
      .dmem_wdata(dmem_wdata),
      .dmem_wstrb(dmem_wstrb),
      .dmem_we   (dmem_we),
      .ebreak    (ebreak)
  );

  //
  // Instruction memory (SRAM)
  //
  svc_mem_sram #(
      .DW       (32),
      .AW       (IMEM_AW),
      .INIT_FILE(IMEM_INIT)
  ) imem (
      .clk    (clk),
      .rst_n  (rst_n),
      .rd_addr(imem_addr),
      .rd_data(imem_data),
      .wr_addr(32'h0),
      .wr_data(32'h0),
      .wr_strb(4'h0),
      .wr_en  (1'b0)
  );

  //
  // Data memory (SRAM)
  //
  svc_mem_sram #(
      .DW(32),
      .AW(DMEM_AW)
  ) dmem (
      .clk    (clk),
      .rst_n  (rst_n),
      .rd_addr(dmem_addr),
      .rd_data(dmem_rdata),
      .wr_addr(dmem_waddr),
      .wr_data(dmem_wdata),
      .wr_strb(dmem_wstrb),
      .wr_en  (dmem_we)
  );

endmodule

`endif
