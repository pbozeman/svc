`ifndef SVC_VGA_MODE_SV
`define SVC_VGA_MODE_SV

// http://www.tinyvga.com/vga-timing/640x480@60Hz
`define VGA_MODE_640x480_H_VISIBLE 640
`define VGA_MODE_640x480_H_FRONT_PORCH 16
`define VGA_MODE_640x480_H_SYNC_PULSE 96
`define VGA_MODE_640x480_H_BACK_PORCH 48
`define VGA_MODE_640x480_H_WHOLE_LINE 800

`define VGA_MODE_640x480_V_VISIBLE 480
`define VGA_MODE_640x480_V_FRONT_PORCH 10
`define VGA_MODE_640x480_V_SYNC_PULSE 2
`define VGA_MODE_640x480_V_BACK_PORCH 33
`define VGA_MODE_640x480_V_WHOLE_FRAME 525

`define VGA_MODE_640x480_H_SYNC_START (`VGA_MODE_640x480_H_VISIBLE + `VGA_MODE_640x480_H_FRONT_PORCH)
`define VGA_MODE_640x480_H_SYNC_END (`VGA_MODE_640x480_H_SYNC_START + `VGA_MODE_640x480_H_SYNC_PULSE)
`define VGA_MODE_640x480_H_LINE_END (`VGA_MODE_640x480_H_WHOLE_LINE - 1)

`define VGA_MODE_640x480_V_SYNC_START (`VGA_MODE_640x480_V_VISIBLE + `VGA_MODE_640x480_V_FRONT_PORCH)
`define VGA_MODE_640x480_V_SYNC_END (`VGA_MODE_640x480_V_SYNC_START + `VGA_MODE_640x480_V_SYNC_PULSE)
`define VGA_MODE_640x480_V_FRAME_END (`VGA_MODE_640x480_V_WHOLE_FRAME - 1)

`endif
