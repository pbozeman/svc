//
// Test case list for svc_cache_axi
//

`TEST_CASE(test_reset);
`TEST_CASE(test_read_miss);
`TEST_CASE(test_read_miss_data);
`TEST_CASE(test_cache_hit);
`TEST_CASE(test_stress);
