`ifndef SVC_VGA_MODE_SV
`define SVC_VGA_MODE_SV

// verilog_format: off

//
// 640x480 60hz
//
// http://www.tinyvga.com/vga-timing/640x480@60Hz
`define VGA_MODE_640x480_H_VISIBLE     640
`define VGA_MODE_640x480_H_FRONT_PORCH 16
`define VGA_MODE_640x480_H_SYNC_PULSE  96
`define VGA_MODE_640x480_H_BACK_PORCH  48
`define VGA_MODE_640x480_H_WHOLE_LINE  800

`define VGA_MODE_640x480_V_VISIBLE     480
`define VGA_MODE_640x480_V_FRONT_PORCH 10
`define VGA_MODE_640x480_V_SYNC_PULSE  2
`define VGA_MODE_640x480_V_BACK_PORCH  33
`define VGA_MODE_640x480_V_WHOLE_FRAME 525

`define VGA_MODE_640x480_H_SYNC_START (`VGA_MODE_640x480_H_VISIBLE    + `VGA_MODE_640x480_H_FRONT_PORCH)
`define VGA_MODE_640x480_H_SYNC_END   (`VGA_MODE_640x480_H_SYNC_START + `VGA_MODE_640x480_H_SYNC_PULSE)
`define VGA_MODE_640x480_H_LINE_END   (`VGA_MODE_640x480_H_WHOLE_LINE - 1)

`define VGA_MODE_640x480_V_SYNC_START (`VGA_MODE_640x480_V_VISIBLE     + `VGA_MODE_640x480_V_FRONT_PORCH)
`define VGA_MODE_640x480_V_SYNC_END   (`VGA_MODE_640x480_V_SYNC_START  + `VGA_MODE_640x480_V_SYNC_PULSE)
`define VGA_MODE_640x480_V_FRAME_END  (`VGA_MODE_640x480_V_WHOLE_FRAME - 1)

`define VGA_MODE_640x480_TB_PIXEL_CLK 40

//
// 800x600 60hz
//
// http://www.tinyvga.com/vga-timing/800x600@60Hz
`define VGA_MODE_800x600_H_VISIBLE     800
`define VGA_MODE_800x600_H_FRONT_PORCH 40
`define VGA_MODE_800x600_H_SYNC_PULSE  128
`define VGA_MODE_800x600_H_BACK_PORCH  88
`define VGA_MODE_800x600_H_WHOLE_LINE  1056

`define VGA_MODE_800x600_V_VISIBLE     600
`define VGA_MODE_800x600_V_FRONT_PORCH 1
`define VGA_MODE_800x600_V_SYNC_PULSE  4
`define VGA_MODE_800x600_V_BACK_PORCH  23
`define VGA_MODE_800x600_V_WHOLE_FRAME 628

`define VGA_MODE_800x600_H_SYNC_START (`VGA_MODE_800x600_H_VISIBLE    + `VGA_MODE_800x600_H_FRONT_PORCH)
`define VGA_MODE_800x600_H_SYNC_END   (`VGA_MODE_800x600_H_SYNC_START + `VGA_MODE_800x600_H_SYNC_PULSE)
`define VGA_MODE_800x600_H_LINE_END   (`VGA_MODE_800x600_H_WHOLE_LINE - 1)

`define VGA_MODE_800x600_V_SYNC_START (`VGA_MODE_800x600_V_VISIBLE     + `VGA_MODE_800x600_V_FRONT_PORCH)
`define VGA_MODE_800x600_V_SYNC_END   (`VGA_MODE_800x600_V_SYNC_START  + `VGA_MODE_800x600_V_SYNC_PULSE)
`define VGA_MODE_800x600_V_FRAME_END  (`VGA_MODE_800x600_V_WHOLE_FRAME - 1)

`define VGA_MODE_800x600_TB_PIXEL_CLK 25

//
// 1024x768 @60hz
// http://www.tinyvga.com/vga-timing/1024x768@60Hz
`define VGA_MODE_1024x768_H_VISIBLE      1024
`define VGA_MODE_1024x768_H_FRONT_PORCH  24
`define VGA_MODE_1024x768_H_SYNC_PULSE   136
`define VGA_MODE_1024x768_H_BACK_PORCH   160
`define VGA_MODE_1024x768_H_WHOLE_LINE   1344

`define VGA_MODE_1024x768_V_VISIBLE      768
`define VGA_MODE_1024x768_V_FRONT_PORCH  3
`define VGA_MODE_1024x768_V_SYNC_PULSE   6
`define VGA_MODE_1024x768_V_BACK_PORCH   29
`define VGA_MODE_1024x768_V_WHOLE_FRAME  806

`define VGA_MODE_1024x768_H_SYNC_START (`VGA_MODE_1024x768_H_VISIBLE    + `VGA_MODE_1024x768_H_FRONT_PORCH)
`define VGA_MODE_1024x768_H_SYNC_END   (`VGA_MODE_1024x768_H_SYNC_START + `VGA_MODE_1024x768_H_SYNC_PULSE)
`define VGA_MODE_1024x768_H_LINE_END   (`VGA_MODE_1024x768_H_WHOLE_LINE - 1)

`define VGA_MODE_1024x768_V_SYNC_START (`VGA_MODE_1024x768_V_VISIBLE     + `VGA_MODE_1024x768_V_FRONT_PORCH)
`define VGA_MODE_1024x768_V_SYNC_END   (`VGA_MODE_1024x768_V_SYNC_START  + `VGA_MODE_1024x768_V_SYNC_PULSE)
`define VGA_MODE_1024x768_V_FRAME_END  (`VGA_MODE_1024x768_V_WHOLE_FRAME - 1)

`define VGA_MODE_1024x768_TB_PIXEL_CLK 15.38

// verilog_format: on
`endif
