`ifndef SVC_ICE40_VGA_MODE_SV
`define SVC_ICE40_VGA_MODE_SV

`include "svc_vga_mode.sv"

// icepll -i 100 -o 25
`define VGA_MODE_640x480_PLL_DIVR (4'd0)
`define VGA_MODE_640x480_PLL_DIVF (7'd7)
`define VGA_MODE_640x480_PLL_DIVQ (3'd5)
`define VGA_MODE_640x480_PLL_FILTER_RANGE (3'd5)

// icepll -i 100 -o 40
`define VGA_MODE_800x600_PLL_DIVR (4'd4)
`define VGA_MODE_800x600_PLL_DIVF (7'd31)
`define VGA_MODE_800x600_PLL_DIVQ (3'd4)
`define VGA_MODE_800x600_PLL_FILTER_RANGE (3'd2)

// icepll -i 100 -o 65
`define VGA_MODE_1024x768_PLL_DIVR (4'd4)
`define VGA_MODE_1024x768_PLL_DIVF (7'd51)
`define VGA_MODE_1024x768_PLL_DIVQ (3'd4)
`define VGA_MODE_1024x768_PLL_FILTER_RANGE (3'd2)

// verilog_format: off
`ifdef VGA_MODE_1024_768_60
  `define VGA_MODE_PLL_DIVR         `VGA_MODE_1024x768_PLL_DIVR
  `define VGA_MODE_PLL_DIVF         `VGA_MODE_1024x768_PLL_DIVF
  `define VGA_MODE_PLL_DIVQ         `VGA_MODE_1024x768_PLL_DIVQ
  `define VGA_MODE_PLL_FILTER_RANGE `VGA_MODE_1024x768_PLL_FILTER_RANGE

  `define VGA_MODE_H_VISIBLE        `VGA_MODE_1024x768_H_VISIBLE
  `define VGA_MODE_H_FRONT_PORCH    `VGA_MODE_1024x768_H_FRONT_PORCH
  `define VGA_MODE_H_SYNC_PULSE     `VGA_MODE_1024x768_H_SYNC_PULSE
  `define VGA_MODE_H_BACK_PORCH     `VGA_MODE_1024x768_H_BACK_PORCH
  `define VGA_MODE_H_WHOLE_LINE     `VGA_MODE_1024x768_H_WHOLE_LINE

  `define VGA_MODE_V_VISIBLE        `VGA_MODE_1024x768_V_VISIBLE
  `define VGA_MODE_V_FRONT_PORCH    `VGA_MODE_1024x768_V_FRONT_PORCH
  `define VGA_MODE_V_SYNC_PULSE     `VGA_MODE_1024x768_V_SYNC_PULSE
  `define VGA_MODE_V_BACK_PORCH     `VGA_MODE_1024x768_V_BACK_PORCH
  `define VGA_MODE_V_WHOLE_FRAME    `VGA_MODE_1024x768_V_WHOLE_FRAME
 
  `define VGA_MODE_TB_PIXEL_CLK     `VGA_MODE_1024x768_TB_PIXEL_CLK
`else
`ifdef VGA_MODE_800_600_60
  `define VGA_MODE_PLL_DIVR         `VGA_MODE_800x600_PLL_DIVR
  `define VGA_MODE_PLL_DIVF         `VGA_MODE_800x600_PLL_DIVF
  `define VGA_MODE_PLL_DIVQ         `VGA_MODE_800x600_PLL_DIVQ
  `define VGA_MODE_PLL_FILTER_RANGE `VGA_MODE_800x600_PLL_FILTER_RANGE

  `define VGA_MODE_H_VISIBLE        `VGA_MODE_800x600_H_VISIBLE
  `define VGA_MODE_H_FRONT_PORCH    `VGA_MODE_800x600_H_FRONT_PORCH
  `define VGA_MODE_H_SYNC_PULSE     `VGA_MODE_800x600_H_SYNC_PULSE
  `define VGA_MODE_H_BACK_PORCH     `VGA_MODE_800x600_H_BACK_PORCH
  `define VGA_MODE_H_WHOLE_LINE     `VGA_MODE_800x600_H_WHOLE_LINE

  `define VGA_MODE_V_VISIBLE        `VGA_MODE_800x600_V_VISIBLE
  `define VGA_MODE_V_FRONT_PORCH    `VGA_MODE_800x600_V_FRONT_PORCH
  `define VGA_MODE_V_SYNC_PULSE     `VGA_MODE_800x600_V_SYNC_PULSE
  `define VGA_MODE_V_BACK_PORCH     `VGA_MODE_800x600_V_BACK_PORCH
  `define VGA_MODE_V_WHOLE_FRAME    `VGA_MODE_800x600_V_WHOLE_FRAME

  `define VGA_MODE_TB_PIXEL_CLK     `VGA_MODE_800x600_TB_PIXEL_CLK
`else
`ifdef VGA_MODE_640_480_60
  `define VGA_MODE_PLL_DIVR         `VGA_MODE_640x480_PLL_DIVR
  `define VGA_MODE_PLL_DIVF         `VGA_MODE_640x480_PLL_DIVF
  `define VGA_MODE_PLL_DIVQ         `VGA_MODE_640x480_PLL_DIVQ
  `define VGA_MODE_PLL_FILTER_RANGE `VGA_MODE_640x480_PLL_FILTER_RANGE

  `define VGA_MODE_H_VISIBLE        `VGA_MODE_640x480_H_VISIBLE
  `define VGA_MODE_H_FRONT_PORCH    `VGA_MODE_640x480_H_FRONT_PORCH
  `define VGA_MODE_H_SYNC_PULSE     `VGA_MODE_640x480_H_SYNC_PULSE
  `define VGA_MODE_H_BACK_PORCH     `VGA_MODE_640x480_H_BACK_PORCH
  `define VGA_MODE_H_WHOLE_LINE     `VGA_MODE_640x480_H_WHOLE_LINE

  `define VGA_MODE_V_VISIBLE        `VGA_MODE_640x480_V_VISIBLE
  `define VGA_MODE_V_FRONT_PORCH    `VGA_MODE_640x480_V_FRONT_PORCH
  `define VGA_MODE_V_SYNC_PULSE     `VGA_MODE_640x480_V_SYNC_PULSE
  `define VGA_MODE_V_BACK_PORCH     `VGA_MODE_640x480_V_BACK_PORCH
  `define VGA_MODE_V_WHOLE_FRAME    `VGA_MODE_640x480_V_WHOLE_FRAME

  `define VGA_MODE_TB_PIXEL_CLK     `VGA_MODE_640x480_TB_PIXEL_CLK
`else
  // There's no `error, so this will have to do
  `include "bad or missing VGA_MODE_ define (consider this an error directive)"
`endif
`endif
`endif

`define VGA_MODE_H_SYNC_START (`VGA_MODE_H_VISIBLE    + `VGA_MODE_H_FRONT_PORCH)
`define VGA_MODE_H_SYNC_END   (`VGA_MODE_H_SYNC_START + `VGA_MODE_H_SYNC_PULSE)
`define VGA_MODE_H_LINE_END   (`VGA_MODE_H_WHOLE_LINE - 1)

`define VGA_MODE_V_SYNC_START (`VGA_MODE_V_VISIBLE    + `VGA_MODE_V_FRONT_PORCH)
`define VGA_MODE_V_SYNC_END   (`VGA_MODE_V_SYNC_START + `VGA_MODE_V_SYNC_PULSE)
`define VGA_MODE_V_FRAME_END  (`VGA_MODE_V_WHOLE_FRAME - 1)
// verilog_format: on

`endif
